module a;real x;initial repeat(50)begin $write("%d",$fscanf(1<<31,"%b",x)==(8*x+1)**0.5%2);end endmodule