module a;integer i,j,x,c;initial begin for(i=0;i<50;i=i+1)begin c=$fscanf(32'h80000000,"%b",x);for(j=0;j<=x;j=j+1)begin c=c+(j*(j+1)/2==x); end $write("%d",c-1);end end endmodule