module c;integer c,d;initial begin while($fscanf(1<<31,"%b",d))begin for(c=1;d>0;c=c+1)d=d-c;$write(~|d);end end endmodule