module z;integer a,b,c,d,e,f,g,h,i,j,k,l,z;initial begin z=$fscanf(1<<31,"%d%d%d%d%d%d%d%d%d%d%d%d",a,b,c,d,e,f,g,h,i,j,k,l);d=d-a;e=e-b;f=f-c;g=g-a;h=h-b;i=i-c;j=j-a;k=k-b;l=l-c;$write((g*k*f+j*e*i+d*h*l-j*h*f-d*k*i-g*e*l)/6);end endmodule